.title KiCad schematic
.include "models/C2012X7R2A104K125AE_p.mod"
.include "models/INA188.lib"
XU2 /INP /INN VEE VDD VSS /GAIN1 /GAIN2 /OUT INA188
XU1 VDD 0 C2012X7R2A104K125AE_p
XU4 0 VEE C2012X7R2A104K125AE_p
XU3 0 VSS C2012X7R2A104K125AE_p
R5 /OUT 0 {RLOAD}
V1 VDD 0 {VPOS}
V3 0 VSS {VNEG}
V4 VEE 0 {VREF}
R1 /IN /INN {RHIGH}
R4 /GAIN1 /GAIN2 {RG}
R2 /INN /INP {RMID}
V2 /IN 0 {VIN}
R3 /INP 0 {RLOW}
.end
